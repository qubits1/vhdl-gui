entity();
