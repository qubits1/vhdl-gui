entity sub3();
