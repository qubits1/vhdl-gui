--new vhdl
