entity sub1();
